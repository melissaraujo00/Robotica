��  CCircuit��  CSerializeHack           ��  CPart            ���  CECapacitor��  CValue  �� ��     4700�F(    U���N@s?      �?�F �� 	 CTerminal  �� ��          �����	@          �  �� ��                              �� ��         ��      �=͈�$�?��  CLED_G�  �� ��                 �          �  ��                             ��          ��      �� 	 CResistor
�  pV �d     560        ��@      �?   �  �h �i         �����	@          �  `h ui         �����	@            td �l         ��      ��  CSPDT��  CToggle   x  �         �  h 1i         �����	@          �  �` a         �����	@          �  �p q                �            \ t          ��    ��  CSPST�  �� ��           �  x� y�               @          �  xx y�          �����	@            t� |�     "      ��    ��  CBattery
�  C� k�     4.5V(          @      �? V �  x� y�                @          �  xy                            l� �     '    ��                  ���  CWire  �� �        *�  ��       *�  �h ��        *�  �h �i       *�  x� y�        *�  �p ��        *�  x�       *�  0h ai       *�  xx �y       *�  �` �y        *�  �` �a                   �                         -    +  0    ,   .  2    2  5   0  " " / # 3 # ' / ' ( ( 1  , 1 + .   - " '   (    # 4 5 3 4    %        �$s�        @     +        @            @    "V  (      �8                
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 