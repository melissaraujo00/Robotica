��  CCircuit��  CSerializeHack           ��  CPart              ���  CNPN��  CDummyValue  `�`�    100hFE            Y@      �? hFE �� 	 CTerminal  `�a�         ��τԠ@V�o��?  �  8�M�        
E����?���2T�?  �  `�a�        s�$�1����t$7��    L�h�         ��      �� 	 CResistor��  CValue  ���    100k        j�@      �?k  �  ��        
E����?���2T��  �  ����     
  �w����!@���2T�?    ���        ��      ��  CBattery�  K�s    9V(          "@      �? V �  ����      
  �w����!@D�t$7��  �  ��!        s�$�1��l�t$7�?    t��         ��      ��  �Vd    120         ^@      �?   �  h)i        ��τԠ@��o���  �  �h�i        $��چ�@��o��?    �dl        ��      ��  CLED_G�  �h�i     	  �w����!@��o��?  �  �h�i        $��چ�@��o���    �\�|    !   ��      ��  CSPST��  CToggle  ����     $   �  ����     
  �w����!@��o��?  �  �x��      	  �w����!@��o���    |���    '     ��    �
�  0� 0�     100hFE            Y@      �? hFE �  0p 1�                 �          �  � �                �          �  0� 1�                              � 8�      +    ��      ��     ,     120         ^@      �?   �  0 11                �          �  �0 1                �            , 4     0    ��      ��  K� s�     9V(          "@      �? V �  �� ��               "@          �  �� ��                             t� ��      4    ��      ��  �0 �1                �          �  �0 �1                �            �$ �D     7    ��      #�%�  �P �p       9   �  �l ��              "@          �  �@ �U                 �            |T �l     ;      ��                  ���  CWire  ����      
 >�  ����      
 >�  `�a!       >�  � a!      >�  `ha�       >�  (hai      >�  �9�      >�  ����     
 >�  �h�i      >�  �h�y      	 >�  �� 1�        >�  0� 1�         >�  00 1q        >�  �0 �1       >�  �0 �A        >�  �0 �1       >�  �� ��                      �                             C   E    A   E  F   ?    B   D  G  ! H ! " " G ' ' @ ( H ( + K + ,   , - - J 0 0 K 1 L 1 4 O 4 5 5 I 7 N 7 8 8 L ; ; O < M < F  ' ?  B  A D   C   @  "  ! ( 5 J - I 0 + 8 1 N < M 7 ; 4   2         �$s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 