��  CCircuit��  CSerializeHack           ��  CPart              ���  CLED_G�� 	 CTerminal   !               �          
�  4 I!               �            44        ��      �� 	 CResistor��  CValue  K� k�     120           ^@      �?   
�  p� q�                 �          
�  p� q�                �            l� t�          ��      ��  CBattery�  �� ��     9V(          "@      �? V 
�  �� ��               "@          
�  �� �               �            �� ��          ��      ��  CSPST��  CToggle  � 0�          
�   � �              "@          
�  ,� A�                �            � ,�            ��    ��  K� s�     4.5V(          @      �? V 
�  ��              @�l1R�-'<  
�  �� ��                  �l1R�-'�    t� �         ��      �
�  �8�9              @�l1R�-'�  
�  �8�9        ��    @�l1R�-'<    �,�L    #    ��      ��  �� �     120           ^@      �?   
�  � 	�          ��    @          
�  � 	        ��    @            � �      '    ��      ��  �� ��       )   
�  �� ��                            
�  �� ��         ��    @            �� ��      +      ��                  ���  CWire  p� q�        .�  @� q�       .�  � 	!      .�  � �!       .�  H q!      .�  p� q!       .�  �� �       .�  �� ��        .�  �8�9      .�  ��9       .�  �� ��        .�  �� ��         .�  	9       .�  �8	9      .�  � 	�        .�  �� 	�                     �                             1    3  /    4  6    2  5    0     8 ! : ! # 7 # $ $ < ' = ' ( ( ; + 9 + , , > 0   / 2   1  4  3 6  5  8 #   7 : + 9 ! ( < $ ; > ' , =            �$s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 