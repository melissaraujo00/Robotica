��  CCircuit��  CSerializeHack           ��  CPart              ��� 
 CVoltmeter��  CMeter  �C�     1.92(    �� 	 CTerminal  P�Q�               @          �  P�Q�        Oo��z�@            D�\�         ��      �� 
 CVResistor��  CSlider  x-�    ��  CValue  R(`    0        @@          
    �  $h9i              @ �3����  �  � hi              @ �3���?    `$t        ��      �� 	 CResistor�  �     120   ������]@      �?   �   )!        Oo��z�@�3���?  �  �  � !                 �3����    � $        ��      ��  CLED�  ����               @ �3���?  �  ���        Oo��z�@ �3����    ����       
 ��      ��  CAmmeter
�  s���     21.5(    �  �x��               @ �3���?  �  ����              @ �3����    ����     #   ��      ��  CBattery�  � �� �    4.5V(          @      �? V �  � �� �               @ �3����  �  � �� �                 �3���?    � �� �     (    ��                    ���  CWire  PhQ�       +�  �hQi      +�  P�Q!       +�  � Q!      +�  �h�y       +�  8h�i      +�  � h� i      +�  � h� �       +�  � �� !        +�  �  � !       +�  � �!       +�  ( �!      +�  ����                     �                             ,    .   1  2    7  5   8    6 # 0 # $ $ 8 ( 3 ( ) ) 4 -  1 ,  / 7 . - #  0 3  2 ( ) 5 4   /  6 $    &        �$s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 