��  CCircuit��  CSerializeHack           ��  CPart              ���  CBattery��  CValue  ����    9V         "@      �? V �� 	 CTerminal  ����             "@          �  ����                            ����        ��      �� 	 CResistor
�  � +�     2.2k          0�@      �?k  �  0� 1�                 �          �  0� 1               �            ,� 4�          ��      ��  CNPN��  CDummyValue  XhXh    100hFE            Y@      �? hFE �  XXYm                �          �  0xEy               �          �  X�Y�     
          �            Dl`�         ��      ��  0H0H    100hFE            Y@      �? hFE �  081M      	          �          �  XY               �          �  0d1y      	        �            L8d         ��      �
�  k���    470k         ��A      �?k  �  ����                �          �  ����               �            ����     "    ��      �
�  �F�T    100k        j�@      �?k  �  �X�Y               �          �  �X�Y               �            �T�\    &    ��                    �              �                                                                  "   " # #   & &   '   '   	         �$s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 