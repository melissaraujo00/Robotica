��  CCircuit��  CSerializeHack           ��  CPart              ��� 	 CInverter�� 	 CTerminal  ����                �          
�  ���     
         @            ����          ��    �
�  p�q�      	        Ğ=          
�  p�q�              @            d�|�          ��    ��  CNPN��  CDummyValue  pppp    100hFE            Y@      �? hFE 
�  p`qu         ��Ş=�� =S;  
�  H�]�        �5��Ş=]�e|�t ;  
�  p�q�     	        Ğ=*� �S�    \tx�         ��      �� 	 CResistor��  CValue  �N\    100k        j�@      �?k  
�  `a        ��Ş=�����Z�:  
�  �`�a        � ��Ş=�����Zݺ    �\d        ��      ��  ����    470k         ��A      �?k  
�  �p��         � ��Ş=s�Aܢ;  
�  ����     	        Ğ=s�Aܢ�    ����         ��      ��  CFloatSwitch��  CWaterLevel  �� ��     	 "   
�  �� ��         �$�Ş=          
�  �� �        b    "@            �� ��      %     ��    ��  CLoudSpeaker�  �)�7    8             @      �?   
�  �(�)        �$�Ş=     \�:  
�  �8�9        ��Ş=     \ƺ    �"�>     *      ��                  �?   ��  CBattery�  ����    9V         "@      �? V 
�  ����       b    "@��b���;  
�  ����     	        Ğ=).s�x�;    ����    /    ��      ��  HPHP    100hFE            Y@      �? hFE 
�  H@IU         m&�Ş=pL�t{^ƺ  
�   `5a        ��Ş=�����Zݺ  
�  HlI�      	 �5��Ş=lM�HE�:    4TPl     3    ��      ��  #� C    2.2k          0�@      �?k  
�  H� I�          �$�Ş=���|^ƺ  
�  HI!        m&�Ş=���|^�:    D� L     8    ��                    ���  CWire  �`�q       ;�  �`�a      ;�  ��q�     	 ;�  p�q�      	 ;�  p�q�      	 ;�  p8qa       ;�  p8�9      ;�  p���     	 ;�  H IA       ;�  p�q�      	 ;�  `!a      ;�  � I�       ;�  � �        ;�  � ��       ;�  ���      ;�   � �       ;�  �� �)       ;�  H� ��                     �                                     ?       A   5    @   F  =   <      > % I % & & K * L * + B + / / J 0 C 0 3 D 3 4 F 4 5 5  8 G 8 9 9 D =  <    E >   C B  A + E 0 9 3 @ ?  4 H M I G H % / K & J M * 8 L           �$s�        @     +        @          ���@    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 