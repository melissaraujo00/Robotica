��  CCircuit��  CSerializeHack           ��  CPart    0   0     ��� 
 CBattery9V��  CDummyValue  � �� �    9V            "@      �? V �� 	 CTerminal  � �� �               .�pj���,�  �  � �� �        ������!@ jC��1�    � �� @         ��   �  ��  CLED�  H�I�        �|�}).�Ԑa�Jf�  �  X�Y�              .�Ԑa�Jf;    A�a�         ����    ��  CLED_Y�  ����     
   Ef�w|).�}�]x�,�  �  �	�              .�}�]x�,;    ���         ����    ��  CLED_G�  ����        �e�z|).����A��  �  ����              .����A�;    ����         ����    �� 	 CResistor
�   ` `    680           @�@      �?   �  `%a        9�|).�``` �$�  �  \`qa        �e�z|).�``` �$;    $Y\i           ��8 	  �
�  h`h`    680           @�@      �?   �  X`ma        9�|).����D7H%�  �  �`�a     
   Ef�w|).����D7H%;    lY�i     "      ��8 	  �
�  �`�`    680           @�@      �?   �  �`�a        9�|).�999y� 5;  �  �`a        �|�}).�999y� 5�    �Y�i     &      ��8 	  ��  CSPST��  CToggle  � ��      )  �  � $� 9       ������!@          �  � $� 9        9�|).�            � �$     ,    ����P    ��  �X�m                �          �  ����                             �l��     /    ��      ��  xXym                �          �  x�y�                             ll��     2    ��      ���  CValue  ��    470         `}@      �?   �  �� �                �          �  �$�9               �            ��$     7    ��      �5�  �    470          `}@      �?   �  �                 �          �  $9               �            $     ;    ��      �5�  Ss    470         `}@      �?   �  x� y                �          �  x$y9               �            t|$     ?    ��      ��  Xm                �          �  ��                             l$�     B    ��      (�*�  �� �      D   �  �� ��              "@          �  �� ��                �            �� ��      F      ��    ��  CBattery5�  3![/    9V(          "@      �? V �  hi              "@          �  h4iI                            \t4     K    ��          0   0     ���  CWire  � 8� �       N�  � 8� 9      N�  (�)      N�  X(	)      N�  �	)       N�  @(Y)      N�  X�Y)       N�  � �A�      N�  @�A)       N�   �I�      N�  ���)       N�   `�       N�  �`��      
 N�  ����     
 N�  p`q�       N�  p���      N�  X89      N�  � y�       N�  �� �       N�  �8Y9      N�  8a       N�  � 8�9      N�  X8Ya       N�  �8�a       N�  �8�Y       N�  x8yY       N�  8Y       N�  x���       N�  �y�       N�  h��       N�  hHi�        N�  x� ��       N�  �� ��        N�  x� y�        N�  � �        N�  h� ��       N�  h� i	           0   0     �    0   0         0   0      V   O    X   U   \   S   ^   Y  c    ] " e " # # [ & f & ' ' Z , , P - - d / g / 0 0 j 2 h 2 3 3 k 7 o 7 8 8 g ; q ; < < i ? p ? @ @ h B i B C C l F r F G G a K s K L L m P  , O R Y T S  Q W U  R  W V T Z   Q ' X # \ [   ^ ]  b c a p G q d e _  - f _ " b & 8 / @ 2 < B 3 0 C j m k L l ` o n 7 n ? ` ; s F r K   I         �$s�        @     +        @            @    "V  (      �P                
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 