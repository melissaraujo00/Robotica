��  CCircuit��  CSerializeHack           ��  CPart              ��� 
 CBattery9V��  CDummyValue  HPHP    9V            "@      �? V �� 	 CTerminal  H@IU                 H�  �   @!U              "@H<    T^�         ��   �  ��  CSPST��  CToggle  �h0�        �  ����             "@          �   ��                             ��0�         ����P    �� 	 CResistor
�  H�H�    680           @�@      �?   �  8�M�             "@H�  �  ����            "@H<    L���           ��8 	  ��  CLED�  �L�a            "@����w?;  �  �L�a             "@����w?�    ��L         ����    ��  CLED_G�  xLya             "@          �  �L�a             "@            q�L          ����    ��  CLED_Y�   T!i             "@          �  0T1i             "@            $9T     $    ����                  ���  CWire  H@A       '�   �A        '�  8@!A      '�  8�9A       '�  ����      '�  �`��       '�  x`yi       '�  0hyi      '�  ����      '�  �`��       '�  �`�i       '�  �h!i                    �                             (   *    ,   )  +    0   1   2     . ! ! - $ $ 3 % % /  )  ( +   * -  ! ,   / % .  1  0  3 2 $   	         �$s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 