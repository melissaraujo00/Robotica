��  CCircuit��  CSerializeHack           ��  CPart              ���  CNPN��  CDummyValue  �� ��     100hFE            Y@      �? hFE �� 	 CTerminal  �� ��                 �          �  �� ��                �          �  ��                             �� �         ��      ��  CSPST��  CToggle  �� ��          �  �� ��              "@          �  �� ��                �            �| ��            ��    �� 	 CResistor��  CValue  pn �|     120         ^@      �?   �  �� ��                �          �  `� u�                �            t| ��         ��      ��  CLED_G�  �� ��                 �          �  �� ��                �            �� ��          ��      ��  h� ��     1k        @�@      �?k  �  �� ��                �          �  X� m�                �            l� ��     "    ��      �� 	 CLDR_Lamp��  CFixedValue  +=9    1M          ��.A      �?M  ��  CLamp  �&�N     %   �  %                �          �  <Q                              $<     *    ��      �� 
 CVResistor��  CSlider   � /�      �  �� �     44k          |�@      �?k 
   0 �  � �                 �          �  � �                �            � �      1    ��      ��  CBattery�  C� k�     9V(          "@      �? V �  x� y�               "@          �  x� y                            l� ��      6    ��                    ���  CWire  �        9�  � �        9�  � Y�       9�  �� ��       9�  � a�       9�  �� �       9�  � �        9�  h�i       9�  xhi       9�  Pi        9�  ��i        9�  xyi        9�  �� ��        9�  �� ��        9�  �� ��       9�  x� ��       9�  x� y�                      �                             F   =    D  I    ?   H  >   G    F " " = # < # * : * + + C 1 @ 1 2 2 ; 6 J 6 7 7 E ; * 2 < : # "  ?   @ > 1 B D E C + A  A 7 B   H   G J  I 6   4         �$s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 