��  CCircuit��  CSerializeHack           ��  CPart              ���  CLED_G�� 	 CTerminal  (` )u          �Q�-� @��~��%�?  
�  (� )�                  ��~��%��    t <�        
 ��      ��  CBattery��  CValue  � � � �     4.5V         @      �? V 
�  � � � �               @��~��%��  
�  � � 	�                 ��~��%�?    � � � �         ��      �� 	 CResistor�  c � � �     120           ^@      �?   
�  � � � �          ��gC6@��~��%��  
�  � � � �               @��~��%�?    � � � �          ��      �� 
 CVResistor��  CSlider  � < � d      �  _ I  W     75          @@033333�?  
    
�  � 0 � E          �Q�-� @��~��%��  
�  � \ � q         ��gC6@��~��%�?    � D � \          ��                    ���  CWire  � � � �        �  � p � �         �  � � � �         �  (� )�          �  � )�         �  (0 )a         �  � 0 )1                     �                             &    $  !    %  "    #  '    " #     !  %  $ '   &            �$s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 